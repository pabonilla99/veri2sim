module not_gate ( input  a, output b );
    assign b = ~a;  // not gate
endmodule
