module and_gate (
    input  a,
    input  b,
    output c
);

    // always @(a or b) begin
    //     c = a & b;
    // end

endmodule
